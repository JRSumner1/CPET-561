
module nios_system (
	clk_clk,
	key_export_export,
	leds_export_export);	

	input		clk_clk;
	input		key_export_export;
	output	[7:0]	leds_export_export;
endmodule
