
module nios_system (
	clk_clk,
	leds_export_export,
	key_export_export);	

	input		clk_clk;
	output	[7:0]	leds_export_export;
	input		key_export_export;
endmodule
